--- !ruby/object:GameState
word:
- E
- u
- r
- i
- p
- i
- d
- e
- a
- n
guessed:
- E
- _
- r
- i
- _
- i
- _
- e
- _
- _
tries: 10
tried_letters:
- e
- l
- m
- i
- r
